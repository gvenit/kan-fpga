    .WEIGHT_CHANNELS(WEIGHT_CHANNELS),