`resetall
`timescale 1ns/1ps
`default_nettype none

/* 
 * MCUWrapperBram : Wrapper for Memory Control Unit
 * 
 * MemoryControlUnit : A Memory Controller that coordinates
 *      the streaming processes for all data, grid and scale 
 *      streams for the data processor.
 * 
 *    The module consists of a global FSM and one local FSM
 *      per output stream. Each FSM may operate with different
 *      clock drivers. The global FSM is expected to work with
 *      the slowest clock of the module.
 * 
 */

module MCUWrapperBram #(
  `include "header_MCUGlobalFSMParameters.vh"
  // BRAM control has ack signal
  parameter BRAM_ACK_SIG = 1,
  // Number of batches per run
  parameter BATCH_SIZE = 1,
  // Width of AXI stream Input Data & Grid interfaces in bits
  parameter DATA_WIDTH = 16,
  // Width of AXI stream Scale interface in bits
  parameter SCALE_WIDTH = 16,
  // Propagate tid signal
  parameter ID_ENABLE = 0,
  // tid signal width
  parameter ID_WIDTH = (ID_ENABLE) ? 8 : 1,
  // Propagate tdest signal
  parameter DEST_ENABLE = 0,
  // tdest signal width
  parameter DEST_WIDTH = (DEST_ENABLE) ? 8 : 1,
  // Propagate tuser signal
  parameter USER_ENABLE = 0,
  // tuser signal width
  parameter USER_WIDTH = (USER_ENABLE) ? 8 : 1,
  // Number of Independent AXI-Stream Data Channels per Batch
  parameter DATA_CHANNELS = 1,
  // Use Common Share Channel 
  parameter SCALE_SHARE = 1,
  // Input Scale Channels
  parameter SCALE_CHANNELS_IN = (SCALE_SHARE)? 1 : DATA_CHANNELS,
  // Output Scale Channels
  parameter SCALE_CHANNELS_OUT = (SCALE_SHARE)? 1 : DATA_CHANNELS*BATCH_SIZE,
  // Use Common Grid Channel 
  parameter GRID_SHARE = 0,
  // Input Grid Channels
  parameter GRID_CHANNELS_IN = (GRID_SHARE)? 1 : DATA_CHANNELS,
  // Output Grid Channels
  parameter GRID_CHANNELS_OUT = (GRID_SHARE)? 1 : DATA_CHANNELS*BATCH_SIZE,
  // Data Width of address bus in bits
  parameter DATA_ADDR = 32,
  // Grid Width of address bus in bits
  parameter GRID_ADDR = 32,
  // Scale Width of address bus in bits
  parameter SCALE_ADDR = 32,
  // Data FIFO size per stream
  parameter DATA_FIFO_DEPTH = (BATCH_SIZE + DATA_CHANNELS),
  // Grid FIFO size per stream
  parameter GRID_FIFO_DEPTH = (BATCH_SIZE + DATA_CHANNELS),
  // Scale FIFO size per stream
  parameter SCALE_FIFO_DEPTH = (SCALE_SHARE) ? 0 : (BATCH_SIZE + DATA_CHANNELS)
) (
  input  wire                                                     fsm_clk,
  input  wire                                                     rst,

  /*
   * Control signals -- Corresponding clock : fsm_clk
   */
  input  wire                                                     operation_start,
  input  wire [DATA_ADDR:0]                                       data_size,
  input  wire [GRID_ADDR:0]                                       grid_size,
  input  wire [SCALE_ADDR:0]                                      scle_size,
  
  /*
   * Interrupt signals -- Corresponding clock : fsm_clk
   */
  output wire                                                     operation_busy,
  output wire                                                     operation_complete,
  output wire                                                     operation_error,

  /*
   * Data BRAM Control Interface -- Corresponding clock : data_bram_clk
   */
  input  wire [BATCH_SIZE*DATA_CHANNELS-1:0]                      data_bram_clk,
  output wire [BATCH_SIZE*DATA_CHANNELS-1:0]                      data_bram_en,
  output wire [BATCH_SIZE*DATA_CHANNELS*DATA_ADDR-1:0]            data_bram_addr,
  input  wire [BATCH_SIZE*DATA_CHANNELS*DATA_WIDTH-1:0]           data_bram_rddata,
  input  wire [BATCH_SIZE*DATA_CHANNELS-1:0]                      data_bram_rdack,  // Ignore if BRAM_ACK_SIG == 0

  /*
   * AXI Stream Data Output -- Corresponding clock : m_axis_data_aclk
   */
  output wire [BATCH_SIZE*DATA_CHANNELS-1:0]                      m_axis_data_aclk,
  output wire [BATCH_SIZE*DATA_CHANNELS*DATA_WIDTH-1:0]           m_axis_data_tdata,
  output wire [BATCH_SIZE*DATA_CHANNELS-1:0]                      m_axis_data_tvalid,
  input  wire [BATCH_SIZE*DATA_CHANNELS-1:0]                      m_axis_data_tready,
  output wire [BATCH_SIZE*DATA_CHANNELS-1:0]                      m_axis_data_tlast,
  output wire [BATCH_SIZE*DATA_CHANNELS*ID_WIDTH-1:0]             m_axis_data_tid,
  output wire [BATCH_SIZE*DATA_CHANNELS*DEST_WIDTH-1:0]           m_axis_data_tdest,
  output wire [BATCH_SIZE*DATA_CHANNELS*USER_WIDTH-1:0]           m_axis_data_tuser,

  /*
   * Grid BRAM Control Interface -- Corresponding clock : grid_bram_clk
   */
  input  wire [GRID_CHANNELS_IN-1:0]                              grid_bram_clk,
  output wire [GRID_CHANNELS_IN-1:0]                              grid_bram_en,
  output wire [GRID_CHANNELS_IN*DATA_ADDR-1:0]                    grid_bram_addr,
  input  wire [GRID_CHANNELS_IN*DATA_WIDTH-1:0]                   grid_bram_rddata,
  input  wire [GRID_CHANNELS_IN-1:0]                              grid_bram_rdack,  // Ignore if BRAM_ACK_SIG == 0                                     

  /*
   * AXI Stream Grid Output -- Corresponding clock : m_axis_grid_aclk
   */
  output wire [GRID_CHANNELS_OUT-1:0]                             m_axis_grid_aclk,
  output wire [GRID_CHANNELS_OUT*DATA_WIDTH-1:0]                  m_axis_grid_tdata,
  output wire [GRID_CHANNELS_OUT-1:0]                             m_axis_grid_tvalid,
  input  wire [GRID_CHANNELS_OUT-1:0]                             m_axis_grid_tready,
  output wire [GRID_CHANNELS_OUT-1:0]                             m_axis_grid_tlast,
  output wire [GRID_CHANNELS_OUT*ID_WIDTH-1:0]                    m_axis_grid_tid,
  output wire [GRID_CHANNELS_OUT*DEST_WIDTH-1:0]                  m_axis_grid_tdest,
  output wire [GRID_CHANNELS_OUT*USER_WIDTH-1:0]                  m_axis_grid_tuser,

  /*
   * Scale BRAM Control Interface -- Corresponding clock : scle_bram_clk
   */
  input  wire [SCALE_CHANNELS_IN-1:0]                             scle_bram_clk,
  output wire [SCALE_CHANNELS_IN-1:0]                             scle_bram_en,
  output wire [SCALE_CHANNELS_IN*SCALE_ADDR-1:0]                  scle_bram_addr,
  input  wire [SCALE_CHANNELS_IN*SCALE_WIDTH-1:0]                 scle_bram_rddata,
  input  wire [SCALE_CHANNELS_IN-1:0]                             scle_bram_rdack,  // Ignore if BRAM_ACK_SIG == 0

  /*
   * AXI Stream Scale Output -- Corresponding clock : m_axis_scle_aclk
   */
  output wire [SCALE_CHANNELS_OUT-1:0]                            m_axis_scle_aclk,
  output wire [SCALE_CHANNELS_OUT*SCALE_WIDTH-1:0]                m_axis_scle_tdata,
  output wire [SCALE_CHANNELS_OUT-1:0]                            m_axis_scle_tvalid,
  input  wire [SCALE_CHANNELS_OUT-1:0]                            m_axis_scle_tready,
  output wire [SCALE_CHANNELS_OUT-1:0]                            m_axis_scle_tlast,
  output wire [SCALE_CHANNELS_OUT*ID_WIDTH-1:0]                   m_axis_scle_tid,
  output wire [SCALE_CHANNELS_OUT*DEST_WIDTH-1:0]                 m_axis_scle_tdest,
  output wire [SCALE_CHANNELS_OUT*USER_WIDTH-1:0]                 m_axis_scle_tuser
);

 MemoryControlUnit #(
  `include "header_MCUGlobalFSMParametersInst.vh"
  // BRAM control has valid signal
  .BRAM_ACK_SIG(BRAM_ACK_SIG),
  // Number of batches per run
  .BATCH_SIZE(BATCH_SIZE),
  // Width of AXI stream Input Data & Grid interfaces in bits
  .DATA_WIDTH(DATA_WIDTH),
  // Width of AXI stream Scale interface in bits
  .SCALE_WIDTH(SCALE_WIDTH),
  // Propagate tid signal
  .ID_ENABLE(ID_ENABLE),
  // tid signal width
  .ID_WIDTH(ID_WIDTH),
  // Propagate tdest signal
  .DEST_ENABLE(DEST_ENABLE),
  // tdest signal width
  .DEST_WIDTH(DEST_WIDTH),
  // Propagate tuser signal
  .USER_ENABLE(USER_ENABLE),
  // tuser signal width
  .USER_WIDTH(USER_WIDTH),
  // Number of Independent AXI-Stream Data Channels per Batch
  .DATA_CHANNELS(DATA_CHANNELS),
  // Use Common Share Channel 
  .SCALE_SHARE(SCALE_SHARE),
  // Input Scale Channels
  .SCALE_CHANNELS_IN(SCALE_CHANNELS_IN),
  // Output Scale Channels
  .SCALE_CHANNELS_OUT(SCALE_CHANNELS_OUT),
  // Use Common Grid Channel 
  .GRID_SHARE(GRID_SHARE),
  // Input Grid Channels
  .GRID_CHANNELS_IN(GRID_CHANNELS_IN),
  // Output Grid Channels
  .GRID_CHANNELS_OUT(GRID_CHANNELS_OUT),
  // Data Width of address bus in bits
  .DATA_ADDR(DATA_ADDR),
  // Grid Width of address bus in bits
  .GRID_ADDR(GRID_ADDR),
  // Scale Width of address bus in bits
  .SCALE_ADDR(SCALE_ADDR),
  // Data FIFO size per stream
  .DATA_FIFO_DEPTH(DATA_FIFO_DEPTH),
  // Grid FIFO size per stream
  .GRID_FIFO_DEPTH(GRID_FIFO_DEPTH),
  // Scale FIFO size per stream
  .SCALE_FIFO_DEPTH(SCALE_FIFO_DEPTH)
 ) mcu_inst (
  .fsm_clk(fsm_clk),
  .rst(rst),
  .operation_start(operation_start),
  .data_size(data_size),
  .grid_size(grid_size),
  .scle_size(scle_size),
  .operation_busy(operation_busy),
  .operation_complete(operation_complete),
  .operation_error(operation_error),
  .data_bram_clk(data_bram_clk),
  .data_bram_en(data_bram_en),
  // .data_bram_we(data_bram_we),
  .data_bram_addr(data_bram_addr),
  // .data_bram_wrdata(data_bram_wrdata),
  .data_bram_rddata(data_bram_rddata),
  .data_bram_rdack(data_bram_rdack),
  .m_axis_data_aclk(m_axis_data_aclk),
  .m_axis_data_tdata(m_axis_data_tdata),
  .m_axis_data_tvalid(m_axis_data_tvalid),
  .m_axis_data_tready(m_axis_data_tready),
  .m_axis_data_tlast(m_axis_data_tlast),
  .m_axis_data_tid(m_axis_data_tid),
  .m_axis_data_tdest(m_axis_data_tdest),
  .m_axis_data_tuser(m_axis_data_tuser),
  .grid_bram_clk(grid_bram_clk),
  .grid_bram_en(grid_bram_en),
  // .grid_bram_we(grid_bram_we),
  .grid_bram_addr(grid_bram_addr),
  // .grid_bram_wrdata(grid_bram_wrdata),
  .grid_bram_rddata(grid_bram_rddata),
  .grid_bram_rdack(grid_bram_rdack),
  .m_axis_grid_aclk(m_axis_grid_aclk),
  .m_axis_grid_tdata(m_axis_grid_tdata),
  .m_axis_grid_tvalid(m_axis_grid_tvalid),
  .m_axis_grid_tready(m_axis_grid_tready),
  .m_axis_grid_tlast(m_axis_grid_tlast),
  .m_axis_grid_tid(m_axis_grid_tid),
  .m_axis_grid_tdest(m_axis_grid_tdest),
  .m_axis_grid_tuser(m_axis_grid_tuser),
  .scle_bram_clk(scle_bram_clk),
  .scle_bram_en(scle_bram_en),
  // .scle_bram_we(scle_bram_we),
  .scle_bram_addr(scle_bram_addr),
  // .scle_bram_wrdata(scle_bram_wrdata),
  .scle_bram_rddata(scle_bram_rddata),
  .scle_bram_rdack(scle_bram_rdack),
  .m_axis_scle_aclk(m_axis_scle_aclk),
  .m_axis_scle_tdata(m_axis_scle_tdata),
  .m_axis_scle_tvalid(m_axis_scle_tvalid),
  .m_axis_scle_tready(m_axis_scle_tready),
  .m_axis_scle_tlast(m_axis_scle_tlast),
  .m_axis_scle_tid(m_axis_scle_tid),
  .m_axis_scle_tdest(m_axis_scle_tdest),
  .m_axis_scle_tuser(m_axis_scle_tuser)
);

endmodule

`resetall
