  parameter NUM_PERIPHERALS = 4,

  // Memory Control Unit
  parameter PERIPHERAL_MCU = 0,
  // Data Processing Unit
  parameter PERIPHERAL_DPU = 1,
  // Axi-Stream Packet Splitter
  parameter PERIPHERAL_APS = 2,
