`ifndef SYSTEM_SIZES_H
`define SYSTEM_SIZES_H
  // Number of Independent AXI-Stream Weight Channels
  parameter WEIGHT_CHANNELS = RSLT_CHANNELS * DATA_CHANNELS,

`endif