    .WEIGHT_CHANNELS(WEIGHT_CHANNELS),
    .GRID_SHARE(GRID_SHARE),
    .SCALE_SHARE(SCALE_SHARE),
    .DATA_CHANNELS_IN(DATA_CHANNELS_IN),
    .DATA_CHANNELS_OUT(DATA_CHANNELS_OUT),
    .RSLT_CHANNELS_OUT(RSLT_CHANNELS_OUT),
    .GRID_CHANNELS_OUT(GRID_CHANNELS_OUT),
    .SCALE_CHANNELS_OUT(SCALE_CHANNELS_OUT),