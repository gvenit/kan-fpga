
  // Global FSM states
  .GLO_FSM_WIDTH(GLO_FSM_WIDTH),
  .GLO_FSM_ST0(GLO_FSM_ST0),
  .GLO_FSM_STR(GLO_FSM_STR),
  .GLO_FSM_OPE(GLO_FSM_OPE),
  .GLO_FSM_END(GLO_FSM_END),
  .GLO_FSM_ERR(GLO_FSM_ERR),
