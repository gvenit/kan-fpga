
  // Global FSM states
  parameter GLO_FSM_WIDTH = 3,
  parameter GLO_FSM_ST0 = 0,
  parameter GLO_FSM_STR = 1,
  parameter GLO_FSM_OPE = 2,
  parameter GLO_FSM_END = 3,
  parameter GLO_FSM_ERR = 4,
